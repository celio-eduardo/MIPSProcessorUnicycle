library verilog;
use verilog.vl_types.all;
entity PCBranch_vlg_vec_tst is
end PCBranch_vlg_vec_tst;
