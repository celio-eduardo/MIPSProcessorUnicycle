library verilog;
use verilog.vl_types.all;
entity JumpEndereco_test_vlg_vec_tst is
end JumpEndereco_test_vlg_vec_tst;
