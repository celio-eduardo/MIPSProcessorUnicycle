library verilog;
use verilog.vl_types.all;
entity mult_divide_vlg_vec_tst is
end mult_divide_vlg_vec_tst;
