library verilog;
use verilog.vl_types.all;
entity DataRamtest_vlg_vec_tst is
end DataRamtest_vlg_vec_tst;
