library verilog;
use verilog.vl_types.all;
entity Controle_ULA_test_vlg_vec_tst is
end Controle_ULA_test_vlg_vec_tst;
